`timescale 1ns / 1ps

module cnn_top #(
    parameter IMG_SIZE = 28,
    parameter DATA_WIDTH = 16,
    parameter CONV1_OUT_CHANNELS = 2,
    parameter CONV2_OUT_CHANNELS = 3,
    parameter CONV1_KERNEL = 5,
    parameter CONV2_KERNEL = 3
)(
    input wire clk,
    input wire reset_n,
    input wire start,
    input wire img_wren,     // Write enable for image RAM
    input wire [9:0]  img_addr,   // <-- expose this pin
	input wire [DATA_WIDTH-1:0]  img_data_in,  // Data to write (if uploading image from host)
    output reg finish,
    output reg [3:0] class_out
);
	// ------------ memory depths -------------
	localparam CONV1_OUT_SIZE = 24;
	localparam MAXRELU1_OUT_SIZE = 12;
	localparam CONV2_OUT_SIZE = 10;
	localparam MAXRELU2_OUT_SIZE = 5;
	localparam FC_OUT_SIZE = 10;
	localparam IMG_PIXELS      = IMG_SIZE*IMG_SIZE; // 784
	localparam W1_WORDS        = CONV1_OUT_CHANNELS*CONV1_KERNEL*CONV1_KERNEL; // 50
	localparam B1_WORDS        = CONV1_OUT_CHANNELS; // 2
	localparam W2_WORDS        = CONV2_OUT_CHANNELS*CONV1_OUT_CHANNELS*CONV2_KERNEL*CONV2_KERNEL; // 54
	localparam B2_WORDS        = CONV2_OUT_CHANNELS; // 3
	localparam WFC_WORDS       = CONV2_OUT_CHANNELS*CONV1_KERNEL*CONV1_KERNEL*CONV2_OUT_SIZE;// 750 
	localparam BFC_WORDS       = FC_OUT_SIZE; // 10
	
	
    // === Wires ===
    (* ramstyle="M4K" *) wire signed [DATA_WIDTH - 1 : 0] conv1_out;
	  wire conv1_finish;
	   
	  (* ramstyle="M4K" *) wire signed [DATA_WIDTH - 1 : 0] max1_out;
	  wire max1_finish;
	 
    (* ramstyle="M4K" *) wire signed [DATA_WIDTH - 1 : 0] conv2_out;
	  wire conv2_finish;
	 
	  (* ramstyle="M4K" *) wire signed [DATA_WIDTH - 1 : 0] max2_out;
	  wire max2_finish;
	 
    (* ramstyle="M4K" *) wire signed [DATA_WIDTH - 1 : 0] fc_out;
	  wire fc_finish;
	 
	  wire argmax_finish;
    
    // Registers for addresses
	reg [9:0] img_addr_counter;       // For image RAM (up to 784 for 28x28)
	reg [5:0] conv1_weight_addr_counter; // For conv1 weights ROM (up to 50)
	reg [0:0] conv1_bias_addr_counter;   // For conv1 bias ROM (up to 2)
	reg [5:0] conv2_weight_addr_counter; // For conv2 weights ROM (up to 54)
	reg [1:0] conv2_bias_addr_counter;   // For conv2 bias ROM (up to 3)
	reg [9:0] fc_weight_addr_counter;  // For fc weights ROM (up to 750) 
    reg [3:0] fc_bias_addr_counter;  // For fc bias ROM (up to 10)
    
    reg [3:0] state;
    wire [3:0] class_predict;
    
    // === FSM VARS ===
    localparam 	S_IDLE 		= 4'd0,
				S_CONV1 	= 4'd1,
				S_MAX1 	 	= 4'd2,
				S_CONV2 	= 4'd3,
				S_MAX2 	 	= 4'd4,
				S_FC 		= 4'd5,
				S_ARGMAX 	= 4'd6,
				S_FINISH 	= 4'd7;
    // === ROMs and RAMs ===
    // Write-side signals (host loads image only while state==S_IDLE)
	// ------------------------------------------------------------------
	wire        wr_en   = (state == S_IDLE) ? img_wren : 1'b0;
	wire [9:0]  wr_addr = (state == S_IDLE) ? img_addr : 10'd0;   // any value when not writing
	wire [DATA_WIDTH-1:0] wr_data = (state == S_IDLE) ? img_data_in : 16'd0;
	
	// Read-side address generated by CNN when running
	// ------------------------------------------------------------------
	wire [9:0]  rd_addr = img_addr_counter;   // your pixel counter
	wire [DATA_WIDTH-1:0] img_data_out;
	// Instantiation of the 2-port, single-clock memory
	// ------------------------------------------------------------------
	img_ram u_img_ram (
		.data      (wr_data),   // 32-bit input
		.wraddress (wr_addr),
		.wren      (wr_en),
		.rdaddress (rd_addr),
		.clock     (clk),       // same clock for both ports
		.q         (img_data_out)
	);
    
	wire [DATA_WIDTH-1:0] conv1_weight_data;

	weight_conv1 rom_conv1_weight (
		.address(conv1_weight_addr_counter),
		.clock(clk),
		.q(conv1_weight_data)
	);
	
	wire [DATA_WIDTH-1:0] conv1_bias_data;

	bias_conv1 rom_conv1_bias (
		.address(conv1_bias_addr_counter),
		.clock(clk),
		.q(conv1_bias_data)
	);
    
	wire [DATA_WIDTH-1:0] conv2_weight_data;

	weight_conv2 rom_conv2_weight (
		.address(conv2_weight_addr_counter),
		.clock(clk),
		.q(conv2_weight_data)
	);
    
	wire [DATA_WIDTH-1:0] conv2_bias_data;

	bias_conv2 rom_conv2_bias (
		.address(conv2_bias_addr_counter),
		.clock(clk),
		.q(conv2_bias_data)
	);
    
	wire [DATA_WIDTH-1:0] fc_weight_data;

	weight_fc rom_fc_weight (
		.address(fc_weight_addr_counter),
		.clock(clk),
		.q(fc_weight_data)
	);
    
	wire [DATA_WIDTH-1:0] fc_bias_data;

	bias_fc rom_fc_bias (
		.address(fc_bias_addr_counter),
		.clock(clk),
		.q(fc_bias_data)
	);
							
		// === Data validation signals ===
		wire data_valid_conv1 = (state == S_CONV1);
		wire result_valid_conv1;
		wire result_valid_max1;
		wire result_valid_conv2;
		wire result_valid_max2;
		wire result_valid_fc;
		integer i;
    
		// === Instantiate modules ===
		wire start_conv1  = (state == S_CONV1);
		wire start_max1   = (state == S_MAX1);
		wire start_conv2  = (state == S_CONV2);
		wire start_max2   = (state == S_MAX2);
		wire start_fc     = (state == S_FC);
		wire start_argmax = (state == S_ARGMAX);
		
		// === Module instances ===
    conv_layer_1 cv1 (
        .clk(clk),
        .reset_n(reset_n),
        .start_conv1(start_conv1),
        .data_valid(data_valid_conv1),
        .partial_image_in(img_data_out),
        .partial_weights_in(conv1_weight_data),
        .partial_biases_in(conv1_bias_data),
        .finish_conv1(conv1_finish),
        .map(conv1_out),
        .result_valid(result_valid_conv1)
    );
    
    maxpool_layer_1 max1 (
        .clk(clk),
        .reset_n(reset_n),
        .start_max1(start_max1),
        .data_valid(result_valid_conv1),
        .data_in(conv1_out),
        .finish_max1(max1_finish),
        .result_valid(result_valid_max1),
        .data_out(max1_out)
    );
    
    conv_layer_2 cv2 (
        .clk(clk),
        .reset_n(reset_n),
        .start_conv2(start_conv2),
        .data_valid(result_valid_max1),
        .partial_image_in(max1_out),
        .partial_weights_in(conv2_weight_data),
        .partial_biases_in(conv2_bias_data),
        .finish_conv2(conv2_finish),
        .map(conv2_out),
        .result_valid(result_valid_conv2)
    );
    
    maxpool_layer_2 max2 (
        .clk(clk),
        .reset_n(reset_n),
        .start_max2(start_max2),
        .data_valid(result_valid_conv2),
        .data_in(conv2_out),
        .finish_max2(max2_finish),
        .result_valid(result_valid_max2),
        .data_out(max2_out)
    );
    
    fc_layer fc (
			.clk(clk),
      .reset_n(reset_n),
      .start_fc(start_fc),
      .data_valid(result_valid_max2),

      // Serial input
      .map_in_serial(max2_out),
      .weight_serial(fc_weight_data),
      .bias_serial(fc_bias_data),

      // Output
      .finish_fc(fc_finish),
      .predict_out(fc_out),
      .predict_out_valid(result_valid_fc)
			);
	 
	 argmax_layer arg (
			.clk(clk),
			.reset_n(reset_n),
			.start_argmax(start_argmax),
			.data_valid(result_valid_fc),
      .class_in(fc_out),
		  .finish_argmax(argmax_finish),
      .index_out(class_predict)
    );
			
			
    
    // === FSM process ===
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            state <= S_IDLE;
            img_addr_counter <= 0;
            conv1_weight_addr_counter <= 0;
            conv1_bias_addr_counter <= 0;
            conv2_weight_addr_counter <= 0;
            conv2_bias_addr_counter <= 0;
            fc_weight_addr_counter <= 0;
            fc_bias_addr_counter <= 0;
            class_out <= 0;
            finish <= 0;
        end else begin
            case (state)
                S_IDLE:     if (start) state <= S_CONV1;
                
                S_CONV1: begin
						if (data_valid_conv1) begin
							if (img_addr_counter < (IMG_PIXELS-1))
								img_addr_counter <= img_addr_counter + 10'b1;
							if (conv1_weight_addr_counter < (W1_WORDS-1))
								conv1_weight_addr_counter <= conv1_weight_addr_counter + 6'b1;
							if (conv1_bias_addr_counter < (B1_WORDS-1))
								conv1_bias_addr_counter <= conv1_bias_addr_counter + 1'b1;
						end
					   if (conv1_finish) state <= S_MAX1;
                end
                
                S_MAX1: begin
					if (max1_finish) state <= S_CONV2;
				end
				
                S_CONV2: begin
						if (result_valid_max1) begin
							if (conv2_weight_addr_counter < (W2_WORDS-1))
								conv2_weight_addr_counter <= conv2_weight_addr_counter + 6'b1;
							if (conv2_bias_addr_counter < (B2_WORDS-1))
								conv2_bias_addr_counter <= conv2_bias_addr_counter + 2'b1;
						end
						if (conv2_finish) state <= S_MAX2;
					end
				
                S_MAX2:     if (max2_finish) state <= S_FC;
                
                S_FC: begin
						if (result_valid_max2) begin
							if (fc_weight_addr_counter < (WFC_WORDS-1))
								fc_weight_addr_counter <= fc_weight_addr_counter + 10'b1;
							if (fc_bias_addr_counter < (BFC_WORDS-1))
								fc_bias_addr_counter <= fc_bias_addr_counter + 4'b1;
						end
						if (fc_finish) state <= S_ARGMAX;
				end
				
				S_ARGMAX:	if (argmax_finish) state <= S_FINISH;
				
                S_FINISH:   begin
					class_out <= class_predict;
					finish <= 1;
					state <= S_IDLE;
                end
                            
                default: begin
					img_addr_counter         <= 0;
					conv1_weight_addr_counter<= 0;
					conv1_bias_addr_counter  <= 0;
					conv2_weight_addr_counter <= 0;
					conv2_bias_addr_counter <= 0;
					fc_weight_addr_counter <= 0;
					fc_bias_addr_counter <= 0;
					state <= S_IDLE;
				end
            endcase
        end
    end
        
endmodule
